//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: router_wrap_tile]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Apr 11 17:54:31 2025
//-------------------------------------------
// ----- BEGIN Grid Verilog module: grid_router_wrap_tile -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for grid_router_wrap_tile -----
module grid_router_wrap_tile(clk_usr,
                             pReset,
                             prog_clk,
                             top_width_0_height_0_subtile_0__pin_data_in_0_,
                             top_width_0_height_0_subtile_0__pin_data_in_1_,
                             top_width_0_height_0_subtile_0__pin_data_in_2_,
                             top_width_0_height_0_subtile_0__pin_data_in_3_,
                             top_width_0_height_0_subtile_0__pin_data_in_4_,
                             top_width_0_height_0_subtile_0__pin_data_in_5_,
                             top_width_0_height_0_subtile_0__pin_data_in_6_,
                             top_width_0_height_0_subtile_0__pin_data_in_7_,
                             top_width_0_height_0_subtile_0__pin_data_in_8_,
                             top_width_0_height_0_subtile_0__pin_data_in_9_,
                             top_width_0_height_0_subtile_0__pin_data_in_10_,
                             top_width_0_height_0_subtile_0__pin_data_in_11_,
                             top_width_0_height_0_subtile_0__pin_data_in_12_,
                             top_width_0_height_0_subtile_0__pin_data_in_13_,
                             top_width_0_height_0_subtile_0__pin_data_in_14_,
                             top_width_0_height_0_subtile_0__pin_data_in_15_,
                             top_width_0_height_0_subtile_0__pin_data_in_16_,
                             top_width_0_height_0_subtile_0__pin_data_in_17_,
                             top_width_0_height_0_subtile_0__pin_data_in_18_,
                             top_width_0_height_0_subtile_0__pin_data_in_19_,
                             top_width_0_height_0_subtile_0__pin_data_in_20_,
                             top_width_0_height_0_subtile_0__pin_data_in_21_,
                             top_width_0_height_0_subtile_0__pin_data_in_22_,
                             top_width_0_height_0_subtile_0__pin_data_in_23_,
                             top_width_0_height_0_subtile_0__pin_data_in_24_,
                             top_width_0_height_0_subtile_0__pin_data_in_25_,
                             top_width_0_height_0_subtile_0__pin_data_in_26_,
                             top_width_0_height_0_subtile_0__pin_data_in_27_,
                             top_width_0_height_0_subtile_0__pin_data_in_28_,
                             top_width_0_height_0_subtile_0__pin_data_in_29_,
                             top_width_0_height_0_subtile_0__pin_data_in_30_,
                             top_width_0_height_0_subtile_0__pin_data_in_31_,
                             top_width_0_height_0_subtile_0__pin_dest_in_0_,
                             top_width_0_height_0_subtile_0__pin_dest_in_1_,
                             top_width_0_height_0_subtile_0__pin_dest_in_2_,
                             top_width_0_height_0_subtile_0__pin_dest_in_3_,
                             top_width_0_height_0_subtile_0__pin_dest_in_4_,
                             top_width_0_height_0_subtile_0__pin_dest_in_5_,
                             top_width_0_height_0_subtile_0__pin_is_tail_in_0_,
                             top_width_0_height_0_subtile_0__pin_send_in_0_,
                             top_width_0_height_0_subtile_0__pin_credit_in_0_,
                             right_width_0_height_1_subtile_0__pin_axis_in_tdest_0_,
                             right_width_0_height_1_subtile_0__pin_axis_in_tdest_1_,
                             right_width_0_height_1_subtile_0__pin_axis_in_tdest_2_,
                             right_width_0_height_1_subtile_0__pin_axis_in_tdest_3_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tready_0_,
                             right_width_0_height_3_subtile_0__pin_data_in_64_,
                             right_width_0_height_3_subtile_0__pin_data_in_65_,
                             right_width_0_height_3_subtile_0__pin_data_in_66_,
                             right_width_0_height_3_subtile_0__pin_data_in_67_,
                             right_width_0_height_3_subtile_0__pin_data_in_68_,
                             right_width_0_height_3_subtile_0__pin_data_in_69_,
                             right_width_0_height_3_subtile_0__pin_data_in_70_,
                             right_width_0_height_3_subtile_0__pin_data_in_71_,
                             right_width_0_height_3_subtile_0__pin_data_in_72_,
                             right_width_0_height_3_subtile_0__pin_data_in_73_,
                             right_width_0_height_3_subtile_0__pin_data_in_74_,
                             right_width_0_height_3_subtile_0__pin_data_in_75_,
                             right_width_0_height_3_subtile_0__pin_data_in_76_,
                             right_width_0_height_3_subtile_0__pin_data_in_77_,
                             right_width_0_height_3_subtile_0__pin_data_in_78_,
                             right_width_0_height_3_subtile_0__pin_data_in_79_,
                             right_width_0_height_3_subtile_0__pin_data_in_80_,
                             right_width_0_height_3_subtile_0__pin_data_in_81_,
                             right_width_0_height_3_subtile_0__pin_data_in_82_,
                             right_width_0_height_3_subtile_0__pin_data_in_83_,
                             right_width_0_height_3_subtile_0__pin_data_in_84_,
                             right_width_0_height_3_subtile_0__pin_data_in_85_,
                             right_width_0_height_3_subtile_0__pin_data_in_86_,
                             right_width_0_height_3_subtile_0__pin_data_in_87_,
                             right_width_0_height_3_subtile_0__pin_data_in_88_,
                             right_width_0_height_3_subtile_0__pin_data_in_89_,
                             right_width_0_height_3_subtile_0__pin_data_in_90_,
                             right_width_0_height_3_subtile_0__pin_data_in_91_,
                             right_width_0_height_3_subtile_0__pin_data_in_92_,
                             right_width_0_height_3_subtile_0__pin_data_in_93_,
                             right_width_0_height_3_subtile_0__pin_data_in_94_,
                             right_width_0_height_3_subtile_0__pin_data_in_95_,
                             right_width_0_height_3_subtile_0__pin_dest_in_6_,
                             right_width_0_height_3_subtile_0__pin_dest_in_7_,
                             right_width_0_height_3_subtile_0__pin_dest_in_8_,
                             right_width_0_height_3_subtile_0__pin_dest_in_9_,
                             right_width_0_height_3_subtile_0__pin_dest_in_10_,
                             right_width_0_height_3_subtile_0__pin_dest_in_11_,
                             right_width_0_height_3_subtile_0__pin_is_tail_in_2_,
                             right_width_0_height_3_subtile_0__pin_send_in_2_,
                             right_width_0_height_3_subtile_0__pin_credit_in_2_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_32_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_33_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_34_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_35_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_36_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_37_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_38_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_39_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_40_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_41_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_42_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_43_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_44_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_45_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_46_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_47_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_48_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_49_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_50_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_51_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_52_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_53_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_54_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_55_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_56_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_57_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_58_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_59_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_60_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_61_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_62_,
                             bottom_width_0_height_0_subtile_0__pin_data_in_63_,
                             bottom_width_0_height_0_subtile_0__pin_dest_in_12_,
                             bottom_width_0_height_0_subtile_0__pin_dest_in_13_,
                             bottom_width_0_height_0_subtile_0__pin_dest_in_14_,
                             bottom_width_0_height_0_subtile_0__pin_dest_in_15_,
                             bottom_width_0_height_0_subtile_0__pin_dest_in_16_,
                             bottom_width_0_height_0_subtile_0__pin_dest_in_17_,
                             bottom_width_0_height_0_subtile_0__pin_is_tail_in_1_,
                             bottom_width_0_height_0_subtile_0__pin_send_in_1_,
                             bottom_width_0_height_0_subtile_0__pin_credit_in_1_,
                             left_width_0_height_0_subtile_0__pin_clk_noc_0_,
                             left_width_0_height_0_subtile_0__pin_rst_n_0_,
                             left_width_0_height_0_subtile_0__pin_router_address_0_,
                             left_width_0_height_0_subtile_0__pin_router_address_1_,
                             left_width_0_height_0_subtile_0__pin_router_address_2_,
                             left_width_0_height_0_subtile_0__pin_router_address_3_,
                             left_width_0_height_0_subtile_0__pin_clk_usr_0_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tvalid_0_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_0_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_1_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_2_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_3_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_4_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_5_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_6_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_7_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_8_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_9_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_10_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_11_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_12_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_13_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_14_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_15_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_16_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_17_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_18_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_19_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_20_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_21_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_22_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_23_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_24_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_25_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_26_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_27_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_28_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_29_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_30_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_31_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_32_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_33_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_34_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_35_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_36_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_37_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_38_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_39_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_40_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_41_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_42_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_43_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_44_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_45_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_46_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_47_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_48_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_49_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_50_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_51_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_52_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_53_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_54_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_55_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_56_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_57_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_58_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_59_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_60_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_61_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_62_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_63_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_64_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_65_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_66_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_67_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_68_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_69_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_70_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_71_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_72_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_73_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_74_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_75_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_76_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_77_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_78_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_79_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_80_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_81_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_82_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_83_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_84_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_85_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_86_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_87_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_88_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_89_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_90_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_91_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_92_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_93_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_94_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_95_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_96_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_97_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_98_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_99_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_100_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_101_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_102_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_103_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_104_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_105_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_106_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_107_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_108_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_109_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_110_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_111_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_112_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_113_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_114_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_115_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_116_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_117_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_118_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_119_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_120_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_121_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_122_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_123_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_124_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_125_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_126_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tdata_127_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tlast_0_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tid_0_,
                             left_width_0_height_1_subtile_0__pin_axis_in_tid_1_,
                             left_width_0_height_3_subtile_0__pin_data_in_96_,
                             left_width_0_height_3_subtile_0__pin_data_in_97_,
                             left_width_0_height_3_subtile_0__pin_data_in_98_,
                             left_width_0_height_3_subtile_0__pin_data_in_99_,
                             left_width_0_height_3_subtile_0__pin_data_in_100_,
                             left_width_0_height_3_subtile_0__pin_data_in_101_,
                             left_width_0_height_3_subtile_0__pin_data_in_102_,
                             left_width_0_height_3_subtile_0__pin_data_in_103_,
                             left_width_0_height_3_subtile_0__pin_data_in_104_,
                             left_width_0_height_3_subtile_0__pin_data_in_105_,
                             left_width_0_height_3_subtile_0__pin_data_in_106_,
                             left_width_0_height_3_subtile_0__pin_data_in_107_,
                             left_width_0_height_3_subtile_0__pin_data_in_108_,
                             left_width_0_height_3_subtile_0__pin_data_in_109_,
                             left_width_0_height_3_subtile_0__pin_data_in_110_,
                             left_width_0_height_3_subtile_0__pin_data_in_111_,
                             left_width_0_height_3_subtile_0__pin_data_in_112_,
                             left_width_0_height_3_subtile_0__pin_data_in_113_,
                             left_width_0_height_3_subtile_0__pin_data_in_114_,
                             left_width_0_height_3_subtile_0__pin_data_in_115_,
                             left_width_0_height_3_subtile_0__pin_data_in_116_,
                             left_width_0_height_3_subtile_0__pin_data_in_117_,
                             left_width_0_height_3_subtile_0__pin_data_in_118_,
                             left_width_0_height_3_subtile_0__pin_data_in_119_,
                             left_width_0_height_3_subtile_0__pin_data_in_120_,
                             left_width_0_height_3_subtile_0__pin_data_in_121_,
                             left_width_0_height_3_subtile_0__pin_data_in_122_,
                             left_width_0_height_3_subtile_0__pin_data_in_123_,
                             left_width_0_height_3_subtile_0__pin_data_in_124_,
                             left_width_0_height_3_subtile_0__pin_data_in_125_,
                             left_width_0_height_3_subtile_0__pin_data_in_126_,
                             left_width_0_height_3_subtile_0__pin_data_in_127_,
                             left_width_0_height_3_subtile_0__pin_dest_in_18_,
                             left_width_0_height_3_subtile_0__pin_dest_in_19_,
                             left_width_0_height_3_subtile_0__pin_dest_in_20_,
                             left_width_0_height_3_subtile_0__pin_dest_in_21_,
                             left_width_0_height_3_subtile_0__pin_dest_in_22_,
                             left_width_0_height_3_subtile_0__pin_dest_in_23_,
                             left_width_0_height_3_subtile_0__pin_is_tail_in_3_,
                             left_width_0_height_3_subtile_0__pin_send_in_3_,
                             left_width_0_height_3_subtile_0__pin_credit_in_3_,
                             ccff_head,
                             top_width_0_height_0_subtile_0__pin_credit_out_0_,
                             top_width_0_height_0_subtile_0__pin_data_out_0_,
                             top_width_0_height_0_subtile_0__pin_data_out_1_,
                             top_width_0_height_0_subtile_0__pin_data_out_2_,
                             top_width_0_height_0_subtile_0__pin_data_out_3_,
                             top_width_0_height_0_subtile_0__pin_data_out_4_,
                             top_width_0_height_0_subtile_0__pin_data_out_5_,
                             top_width_0_height_0_subtile_0__pin_data_out_6_,
                             top_width_0_height_0_subtile_0__pin_data_out_7_,
                             top_width_0_height_0_subtile_0__pin_data_out_8_,
                             top_width_0_height_0_subtile_0__pin_data_out_9_,
                             top_width_0_height_0_subtile_0__pin_data_out_10_,
                             top_width_0_height_0_subtile_0__pin_data_out_11_,
                             top_width_0_height_0_subtile_0__pin_data_out_12_,
                             top_width_0_height_0_subtile_0__pin_data_out_13_,
                             top_width_0_height_0_subtile_0__pin_data_out_14_,
                             top_width_0_height_0_subtile_0__pin_data_out_15_,
                             top_width_0_height_0_subtile_0__pin_data_out_16_,
                             top_width_0_height_0_subtile_0__pin_data_out_17_,
                             top_width_0_height_0_subtile_0__pin_data_out_18_,
                             top_width_0_height_0_subtile_0__pin_data_out_19_,
                             top_width_0_height_0_subtile_0__pin_data_out_20_,
                             top_width_0_height_0_subtile_0__pin_data_out_21_,
                             top_width_0_height_0_subtile_0__pin_data_out_22_,
                             top_width_0_height_0_subtile_0__pin_data_out_23_,
                             top_width_0_height_0_subtile_0__pin_data_out_24_,
                             top_width_0_height_0_subtile_0__pin_data_out_25_,
                             top_width_0_height_0_subtile_0__pin_data_out_26_,
                             top_width_0_height_0_subtile_0__pin_data_out_27_,
                             top_width_0_height_0_subtile_0__pin_data_out_28_,
                             top_width_0_height_0_subtile_0__pin_data_out_29_,
                             top_width_0_height_0_subtile_0__pin_data_out_30_,
                             top_width_0_height_0_subtile_0__pin_data_out_31_,
                             top_width_0_height_0_subtile_0__pin_dest_out_0_,
                             top_width_0_height_0_subtile_0__pin_dest_out_1_,
                             top_width_0_height_0_subtile_0__pin_dest_out_2_,
                             top_width_0_height_0_subtile_0__pin_dest_out_3_,
                             top_width_0_height_0_subtile_0__pin_dest_out_4_,
                             top_width_0_height_0_subtile_0__pin_dest_out_5_,
                             top_width_0_height_0_subtile_0__pin_is_tail_out_0_,
                             top_width_0_height_0_subtile_0__pin_send_out_0_,
                             right_width_0_height_0_subtile_0__pin_axis_in_tready_0_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tlast_0_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tid_0_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tid_1_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tdest_0_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tdest_1_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tdest_2_,
                             right_width_0_height_0_subtile_0__pin_axis_out_tdest_3_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tvalid_0_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_0_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_1_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_2_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_3_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_4_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_5_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_6_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_7_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_8_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_9_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_10_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_11_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_12_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_13_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_14_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_15_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_16_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_17_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_18_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_19_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_20_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_21_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_22_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_23_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_24_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_25_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_26_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_27_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_28_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_29_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_30_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_31_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_32_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_33_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_34_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_35_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_36_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_37_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_38_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_39_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_40_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_41_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_42_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_43_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_44_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_45_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_46_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_47_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_48_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_49_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_50_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_51_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_52_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_53_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_54_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_55_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_56_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_57_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_58_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_59_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_60_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_61_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_62_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_63_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_64_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_65_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_66_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_67_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_68_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_69_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_70_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_71_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_72_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_73_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_74_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_75_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_76_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_77_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_78_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_79_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_80_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_81_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_82_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_83_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_84_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_85_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_86_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_87_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_88_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_89_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_90_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_91_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_92_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_93_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_94_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_95_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_96_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_97_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_98_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_99_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_100_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_101_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_102_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_103_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_104_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_105_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_106_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_107_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_108_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_109_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_110_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_111_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_112_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_113_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_114_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_115_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_116_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_117_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_118_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_119_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_120_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_121_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_122_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_123_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_124_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_125_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_126_,
                             right_width_0_height_1_subtile_0__pin_axis_out_tdata_127_,
                             right_width_0_height_3_subtile_0__pin_credit_out_2_,
                             right_width_0_height_3_subtile_0__pin_data_out_64_,
                             right_width_0_height_3_subtile_0__pin_data_out_65_,
                             right_width_0_height_3_subtile_0__pin_data_out_66_,
                             right_width_0_height_3_subtile_0__pin_data_out_67_,
                             right_width_0_height_3_subtile_0__pin_data_out_68_,
                             right_width_0_height_3_subtile_0__pin_data_out_69_,
                             right_width_0_height_3_subtile_0__pin_data_out_70_,
                             right_width_0_height_3_subtile_0__pin_data_out_71_,
                             right_width_0_height_3_subtile_0__pin_data_out_72_,
                             right_width_0_height_3_subtile_0__pin_data_out_73_,
                             right_width_0_height_3_subtile_0__pin_data_out_74_,
                             right_width_0_height_3_subtile_0__pin_data_out_75_,
                             right_width_0_height_3_subtile_0__pin_data_out_76_,
                             right_width_0_height_3_subtile_0__pin_data_out_77_,
                             right_width_0_height_3_subtile_0__pin_data_out_78_,
                             right_width_0_height_3_subtile_0__pin_data_out_79_,
                             right_width_0_height_3_subtile_0__pin_data_out_80_,
                             right_width_0_height_3_subtile_0__pin_data_out_81_,
                             right_width_0_height_3_subtile_0__pin_data_out_82_,
                             right_width_0_height_3_subtile_0__pin_data_out_83_,
                             right_width_0_height_3_subtile_0__pin_data_out_84_,
                             right_width_0_height_3_subtile_0__pin_data_out_85_,
                             right_width_0_height_3_subtile_0__pin_data_out_86_,
                             right_width_0_height_3_subtile_0__pin_data_out_87_,
                             right_width_0_height_3_subtile_0__pin_data_out_88_,
                             right_width_0_height_3_subtile_0__pin_data_out_89_,
                             right_width_0_height_3_subtile_0__pin_data_out_90_,
                             right_width_0_height_3_subtile_0__pin_data_out_91_,
                             right_width_0_height_3_subtile_0__pin_data_out_92_,
                             right_width_0_height_3_subtile_0__pin_data_out_93_,
                             right_width_0_height_3_subtile_0__pin_data_out_94_,
                             right_width_0_height_3_subtile_0__pin_data_out_95_,
                             right_width_0_height_3_subtile_0__pin_dest_out_6_,
                             right_width_0_height_3_subtile_0__pin_dest_out_7_,
                             right_width_0_height_3_subtile_0__pin_dest_out_8_,
                             right_width_0_height_3_subtile_0__pin_dest_out_9_,
                             right_width_0_height_3_subtile_0__pin_dest_out_10_,
                             right_width_0_height_3_subtile_0__pin_dest_out_11_,
                             right_width_0_height_3_subtile_0__pin_is_tail_out_2_,
                             right_width_0_height_3_subtile_0__pin_send_out_2_,
                             bottom_width_0_height_0_subtile_0__pin_credit_out_1_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_32_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_33_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_34_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_35_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_36_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_37_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_38_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_39_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_40_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_41_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_42_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_43_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_44_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_45_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_46_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_47_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_48_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_49_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_50_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_51_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_52_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_53_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_54_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_55_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_56_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_57_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_58_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_59_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_60_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_61_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_62_,
                             bottom_width_0_height_0_subtile_0__pin_data_out_63_,
                             bottom_width_0_height_0_subtile_0__pin_dest_out_12_,
                             bottom_width_0_height_0_subtile_0__pin_dest_out_13_,
                             bottom_width_0_height_0_subtile_0__pin_dest_out_14_,
                             bottom_width_0_height_0_subtile_0__pin_dest_out_15_,
                             bottom_width_0_height_0_subtile_0__pin_dest_out_16_,
                             bottom_width_0_height_0_subtile_0__pin_dest_out_17_,
                             bottom_width_0_height_0_subtile_0__pin_is_tail_out_1_,
                             bottom_width_0_height_0_subtile_0__pin_send_out_1_,
                             left_width_0_height_3_subtile_0__pin_credit_out_3_,
                             left_width_0_height_3_subtile_0__pin_data_out_96_,
                             left_width_0_height_3_subtile_0__pin_data_out_97_,
                             left_width_0_height_3_subtile_0__pin_data_out_98_,
                             left_width_0_height_3_subtile_0__pin_data_out_99_,
                             left_width_0_height_3_subtile_0__pin_data_out_100_,
                             left_width_0_height_3_subtile_0__pin_data_out_101_,
                             left_width_0_height_3_subtile_0__pin_data_out_102_,
                             left_width_0_height_3_subtile_0__pin_data_out_103_,
                             left_width_0_height_3_subtile_0__pin_data_out_104_,
                             left_width_0_height_3_subtile_0__pin_data_out_105_,
                             left_width_0_height_3_subtile_0__pin_data_out_106_,
                             left_width_0_height_3_subtile_0__pin_data_out_107_,
                             left_width_0_height_3_subtile_0__pin_data_out_108_,
                             left_width_0_height_3_subtile_0__pin_data_out_109_,
                             left_width_0_height_3_subtile_0__pin_data_out_110_,
                             left_width_0_height_3_subtile_0__pin_data_out_111_,
                             left_width_0_height_3_subtile_0__pin_data_out_112_,
                             left_width_0_height_3_subtile_0__pin_data_out_113_,
                             left_width_0_height_3_subtile_0__pin_data_out_114_,
                             left_width_0_height_3_subtile_0__pin_data_out_115_,
                             left_width_0_height_3_subtile_0__pin_data_out_116_,
                             left_width_0_height_3_subtile_0__pin_data_out_117_,
                             left_width_0_height_3_subtile_0__pin_data_out_118_,
                             left_width_0_height_3_subtile_0__pin_data_out_119_,
                             left_width_0_height_3_subtile_0__pin_data_out_120_,
                             left_width_0_height_3_subtile_0__pin_data_out_121_,
                             left_width_0_height_3_subtile_0__pin_data_out_122_,
                             left_width_0_height_3_subtile_0__pin_data_out_123_,
                             left_width_0_height_3_subtile_0__pin_data_out_124_,
                             left_width_0_height_3_subtile_0__pin_data_out_125_,
                             left_width_0_height_3_subtile_0__pin_data_out_126_,
                             left_width_0_height_3_subtile_0__pin_data_out_127_,
                             left_width_0_height_3_subtile_0__pin_dest_out_13_,
                             left_width_0_height_3_subtile_0__pin_dest_out_14_,
                             left_width_0_height_3_subtile_0__pin_dest_out_15_,
                             left_width_0_height_3_subtile_0__pin_dest_out_16_,
                             left_width_0_height_3_subtile_0__pin_dest_out_17_,
                             left_width_0_height_3_subtile_0__pin_dest_out_18_,
                             left_width_0_height_3_subtile_0__pin_dest_out_19_,
                             left_width_0_height_3_subtile_0__pin_dest_out_20_,
                             left_width_0_height_3_subtile_0__pin_dest_out_21_,
                             left_width_0_height_3_subtile_0__pin_dest_out_22_,
                             left_width_0_height_3_subtile_0__pin_dest_out_23_,
                             left_width_0_height_3_subtile_0__pin_is_tail_out_3_,
                             left_width_0_height_3_subtile_0__pin_send_out_3_,
                             ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk_usr;
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_data_in_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_dest_in_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_dest_in_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_dest_in_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_dest_in_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_dest_in_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_dest_in_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_is_tail_in_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_send_in_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_credit_in_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_axis_in_tdest_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_axis_in_tdest_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_axis_in_tdest_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_axis_in_tdest_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tready_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_64_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_65_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_66_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_67_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_68_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_69_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_70_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_71_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_72_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_73_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_74_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_75_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_76_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_77_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_78_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_79_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_80_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_81_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_82_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_83_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_84_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_85_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_86_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_87_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_88_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_89_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_90_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_91_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_92_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_93_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_94_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_data_in_95_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_dest_in_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_dest_in_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_dest_in_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_dest_in_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_dest_in_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_dest_in_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_is_tail_in_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_send_in_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_credit_in_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_32_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_33_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_34_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_35_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_36_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_37_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_38_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_39_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_40_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_41_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_42_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_43_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_44_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_45_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_46_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_47_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_48_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_49_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_50_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_51_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_52_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_53_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_54_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_55_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_56_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_57_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_58_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_59_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_60_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_61_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_62_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_data_in_63_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_dest_in_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_dest_in_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_dest_in_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_dest_in_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_dest_in_16_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_dest_in_17_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_is_tail_in_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_send_in_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_credit_in_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_noc_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_rst_n_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_router_address_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_router_address_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_router_address_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_router_address_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_usr_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tvalid_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_19_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_20_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_21_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_22_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_23_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_24_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_25_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_26_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_27_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_28_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_29_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_30_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_31_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_32_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_33_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_34_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_35_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_36_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_37_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_38_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_39_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_40_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_41_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_42_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_43_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_44_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_45_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_46_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_47_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_48_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_49_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_50_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_51_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_52_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_53_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_54_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_55_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_56_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_57_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_58_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_59_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_60_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_61_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_62_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_63_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_64_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_65_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_66_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_67_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_68_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_69_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_70_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_71_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_72_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_73_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_74_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_75_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_76_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_77_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_78_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_79_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_80_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_81_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_82_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_83_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_84_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_85_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_86_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_87_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_88_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_89_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_90_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_91_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_92_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_93_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_94_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_95_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_96_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_97_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_98_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_99_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_100_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_101_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_102_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_103_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_104_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_105_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_106_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_107_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_108_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_109_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_110_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_111_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_112_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_113_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_114_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_115_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_116_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_117_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_118_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_119_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_120_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_121_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_122_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_123_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_124_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_125_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_126_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tdata_127_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tlast_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tid_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_axis_in_tid_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_96_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_97_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_98_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_99_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_100_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_101_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_102_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_103_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_104_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_105_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_106_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_107_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_108_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_109_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_110_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_111_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_112_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_113_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_114_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_115_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_116_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_117_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_118_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_119_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_120_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_121_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_122_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_123_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_124_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_125_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_126_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_data_in_127_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_dest_in_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_dest_in_19_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_dest_in_20_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_dest_in_21_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_dest_in_22_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_dest_in_23_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_is_tail_in_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_send_in_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_3_subtile_0__pin_credit_in_3_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_credit_out_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_12_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_13_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_14_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_15_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_16_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_17_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_18_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_19_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_20_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_21_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_22_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_23_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_24_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_25_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_26_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_27_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_28_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_29_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_30_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_data_out_31_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_dest_out_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_dest_out_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_dest_out_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_dest_out_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_dest_out_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_dest_out_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_is_tail_out_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_send_out_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_in_tready_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tlast_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tid_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tid_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tdest_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tdest_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tdest_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_axis_out_tdest_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tvalid_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_24_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_25_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_26_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_27_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_28_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_29_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_30_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_31_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_32_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_33_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_34_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_35_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_36_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_37_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_38_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_39_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_40_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_41_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_42_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_43_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_44_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_45_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_46_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_47_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_48_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_49_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_50_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_51_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_52_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_53_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_54_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_55_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_56_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_57_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_58_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_59_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_60_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_61_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_62_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_63_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_64_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_65_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_66_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_67_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_68_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_69_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_70_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_71_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_72_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_73_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_74_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_75_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_76_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_77_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_78_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_79_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_80_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_81_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_82_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_83_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_84_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_85_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_86_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_87_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_88_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_89_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_90_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_91_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_92_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_93_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_94_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_95_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_96_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_97_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_98_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_99_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_100_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_101_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_102_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_103_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_104_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_105_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_106_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_107_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_108_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_109_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_110_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_111_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_112_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_113_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_114_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_115_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_116_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_117_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_118_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_119_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_120_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_121_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_122_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_123_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_124_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_125_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_126_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_axis_out_tdata_127_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_credit_out_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_64_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_65_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_66_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_67_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_68_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_69_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_70_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_71_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_72_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_73_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_74_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_75_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_76_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_77_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_78_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_79_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_80_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_81_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_82_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_83_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_84_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_85_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_86_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_87_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_88_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_89_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_90_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_91_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_92_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_93_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_94_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_data_out_95_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_dest_out_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_dest_out_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_dest_out_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_dest_out_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_dest_out_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_dest_out_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_is_tail_out_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_send_out_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_credit_out_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_33_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_34_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_35_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_36_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_37_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_38_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_39_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_40_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_41_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_42_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_43_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_44_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_45_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_46_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_47_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_48_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_49_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_50_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_51_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_52_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_53_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_54_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_55_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_56_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_57_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_58_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_59_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_60_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_61_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_62_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_data_out_63_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_dest_out_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_dest_out_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_dest_out_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_dest_out_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_dest_out_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_dest_out_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_is_tail_out_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_send_out_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_credit_out_3_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_96_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_97_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_98_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_99_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_100_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_101_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_102_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_103_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_104_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_105_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_106_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_107_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_108_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_109_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_110_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_111_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_112_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_113_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_114_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_115_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_116_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_117_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_118_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_119_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_120_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_121_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_122_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_123_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_124_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_125_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_126_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_data_out_127_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_13_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_14_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_15_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_16_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_17_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_18_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_19_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_20_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_21_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_22_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_dest_out_23_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_is_tail_out_3_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_3_subtile_0__pin_send_out_3_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [13:17] logical_tile_router_wrap_tile_mode_router_wrap_tile__0_undriven_router_wrap_tile_dest_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_router_wrap_tile_mode_router_wrap_tile_ logical_tile_router_wrap_tile_mode_router_wrap_tile__0 (
		.clk_usr(clk_usr),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.router_wrap_tile_clk_noc(left_width_0_height_0_subtile_0__pin_clk_noc_0_),
		.router_wrap_tile_rst_n(left_width_0_height_0_subtile_0__pin_rst_n_0_),
		.router_wrap_tile_data_in({top_width_0_height_0_subtile_0__pin_data_in_0_, top_width_0_height_0_subtile_0__pin_data_in_1_, top_width_0_height_0_subtile_0__pin_data_in_2_, top_width_0_height_0_subtile_0__pin_data_in_3_, top_width_0_height_0_subtile_0__pin_data_in_4_, top_width_0_height_0_subtile_0__pin_data_in_5_, top_width_0_height_0_subtile_0__pin_data_in_6_, top_width_0_height_0_subtile_0__pin_data_in_7_, top_width_0_height_0_subtile_0__pin_data_in_8_, top_width_0_height_0_subtile_0__pin_data_in_9_, top_width_0_height_0_subtile_0__pin_data_in_10_, top_width_0_height_0_subtile_0__pin_data_in_11_, top_width_0_height_0_subtile_0__pin_data_in_12_, top_width_0_height_0_subtile_0__pin_data_in_13_, top_width_0_height_0_subtile_0__pin_data_in_14_, top_width_0_height_0_subtile_0__pin_data_in_15_, top_width_0_height_0_subtile_0__pin_data_in_16_, top_width_0_height_0_subtile_0__pin_data_in_17_, top_width_0_height_0_subtile_0__pin_data_in_18_, top_width_0_height_0_subtile_0__pin_data_in_19_, top_width_0_height_0_subtile_0__pin_data_in_20_, top_width_0_height_0_subtile_0__pin_data_in_21_, top_width_0_height_0_subtile_0__pin_data_in_22_, top_width_0_height_0_subtile_0__pin_data_in_23_, top_width_0_height_0_subtile_0__pin_data_in_24_, top_width_0_height_0_subtile_0__pin_data_in_25_, top_width_0_height_0_subtile_0__pin_data_in_26_, top_width_0_height_0_subtile_0__pin_data_in_27_, top_width_0_height_0_subtile_0__pin_data_in_28_, top_width_0_height_0_subtile_0__pin_data_in_29_, top_width_0_height_0_subtile_0__pin_data_in_30_, top_width_0_height_0_subtile_0__pin_data_in_31_, bottom_width_0_height_0_subtile_0__pin_data_in_32_, bottom_width_0_height_0_subtile_0__pin_data_in_33_, bottom_width_0_height_0_subtile_0__pin_data_in_34_, bottom_width_0_height_0_subtile_0__pin_data_in_35_, bottom_width_0_height_0_subtile_0__pin_data_in_36_, bottom_width_0_height_0_subtile_0__pin_data_in_37_, bottom_width_0_height_0_subtile_0__pin_data_in_38_, bottom_width_0_height_0_subtile_0__pin_data_in_39_, bottom_width_0_height_0_subtile_0__pin_data_in_40_, bottom_width_0_height_0_subtile_0__pin_data_in_41_, bottom_width_0_height_0_subtile_0__pin_data_in_42_, bottom_width_0_height_0_subtile_0__pin_data_in_43_, bottom_width_0_height_0_subtile_0__pin_data_in_44_, bottom_width_0_height_0_subtile_0__pin_data_in_45_, bottom_width_0_height_0_subtile_0__pin_data_in_46_, bottom_width_0_height_0_subtile_0__pin_data_in_47_, bottom_width_0_height_0_subtile_0__pin_data_in_48_, bottom_width_0_height_0_subtile_0__pin_data_in_49_, bottom_width_0_height_0_subtile_0__pin_data_in_50_, bottom_width_0_height_0_subtile_0__pin_data_in_51_, bottom_width_0_height_0_subtile_0__pin_data_in_52_, bottom_width_0_height_0_subtile_0__pin_data_in_53_, bottom_width_0_height_0_subtile_0__pin_data_in_54_, bottom_width_0_height_0_subtile_0__pin_data_in_55_, bottom_width_0_height_0_subtile_0__pin_data_in_56_, bottom_width_0_height_0_subtile_0__pin_data_in_57_, bottom_width_0_height_0_subtile_0__pin_data_in_58_, bottom_width_0_height_0_subtile_0__pin_data_in_59_, bottom_width_0_height_0_subtile_0__pin_data_in_60_, bottom_width_0_height_0_subtile_0__pin_data_in_61_, bottom_width_0_height_0_subtile_0__pin_data_in_62_, bottom_width_0_height_0_subtile_0__pin_data_in_63_, right_width_0_height_3_subtile_0__pin_data_in_64_, right_width_0_height_3_subtile_0__pin_data_in_65_, right_width_0_height_3_subtile_0__pin_data_in_66_, right_width_0_height_3_subtile_0__pin_data_in_67_, right_width_0_height_3_subtile_0__pin_data_in_68_, right_width_0_height_3_subtile_0__pin_data_in_69_, right_width_0_height_3_subtile_0__pin_data_in_70_, right_width_0_height_3_subtile_0__pin_data_in_71_, right_width_0_height_3_subtile_0__pin_data_in_72_, right_width_0_height_3_subtile_0__pin_data_in_73_, right_width_0_height_3_subtile_0__pin_data_in_74_, right_width_0_height_3_subtile_0__pin_data_in_75_, right_width_0_height_3_subtile_0__pin_data_in_76_, right_width_0_height_3_subtile_0__pin_data_in_77_, right_width_0_height_3_subtile_0__pin_data_in_78_, right_width_0_height_3_subtile_0__pin_data_in_79_, right_width_0_height_3_subtile_0__pin_data_in_80_, right_width_0_height_3_subtile_0__pin_data_in_81_, right_width_0_height_3_subtile_0__pin_data_in_82_, right_width_0_height_3_subtile_0__pin_data_in_83_, right_width_0_height_3_subtile_0__pin_data_in_84_, right_width_0_height_3_subtile_0__pin_data_in_85_, right_width_0_height_3_subtile_0__pin_data_in_86_, right_width_0_height_3_subtile_0__pin_data_in_87_, right_width_0_height_3_subtile_0__pin_data_in_88_, right_width_0_height_3_subtile_0__pin_data_in_89_, right_width_0_height_3_subtile_0__pin_data_in_90_, right_width_0_height_3_subtile_0__pin_data_in_91_, right_width_0_height_3_subtile_0__pin_data_in_92_, right_width_0_height_3_subtile_0__pin_data_in_93_, right_width_0_height_3_subtile_0__pin_data_in_94_, right_width_0_height_3_subtile_0__pin_data_in_95_, left_width_0_height_3_subtile_0__pin_data_in_96_, left_width_0_height_3_subtile_0__pin_data_in_97_, left_width_0_height_3_subtile_0__pin_data_in_98_, left_width_0_height_3_subtile_0__pin_data_in_99_, left_width_0_height_3_subtile_0__pin_data_in_100_, left_width_0_height_3_subtile_0__pin_data_in_101_, left_width_0_height_3_subtile_0__pin_data_in_102_, left_width_0_height_3_subtile_0__pin_data_in_103_, left_width_0_height_3_subtile_0__pin_data_in_104_, left_width_0_height_3_subtile_0__pin_data_in_105_, left_width_0_height_3_subtile_0__pin_data_in_106_, left_width_0_height_3_subtile_0__pin_data_in_107_, left_width_0_height_3_subtile_0__pin_data_in_108_, left_width_0_height_3_subtile_0__pin_data_in_109_, left_width_0_height_3_subtile_0__pin_data_in_110_, left_width_0_height_3_subtile_0__pin_data_in_111_, left_width_0_height_3_subtile_0__pin_data_in_112_, left_width_0_height_3_subtile_0__pin_data_in_113_, left_width_0_height_3_subtile_0__pin_data_in_114_, left_width_0_height_3_subtile_0__pin_data_in_115_, left_width_0_height_3_subtile_0__pin_data_in_116_, left_width_0_height_3_subtile_0__pin_data_in_117_, left_width_0_height_3_subtile_0__pin_data_in_118_, left_width_0_height_3_subtile_0__pin_data_in_119_, left_width_0_height_3_subtile_0__pin_data_in_120_, left_width_0_height_3_subtile_0__pin_data_in_121_, left_width_0_height_3_subtile_0__pin_data_in_122_, left_width_0_height_3_subtile_0__pin_data_in_123_, left_width_0_height_3_subtile_0__pin_data_in_124_, left_width_0_height_3_subtile_0__pin_data_in_125_, left_width_0_height_3_subtile_0__pin_data_in_126_, left_width_0_height_3_subtile_0__pin_data_in_127_}),
		.router_wrap_tile_dest_in({top_width_0_height_0_subtile_0__pin_dest_in_0_, top_width_0_height_0_subtile_0__pin_dest_in_1_, top_width_0_height_0_subtile_0__pin_dest_in_2_, top_width_0_height_0_subtile_0__pin_dest_in_3_, top_width_0_height_0_subtile_0__pin_dest_in_4_, top_width_0_height_0_subtile_0__pin_dest_in_5_, right_width_0_height_3_subtile_0__pin_dest_in_6_, right_width_0_height_3_subtile_0__pin_dest_in_7_, right_width_0_height_3_subtile_0__pin_dest_in_8_, right_width_0_height_3_subtile_0__pin_dest_in_9_, right_width_0_height_3_subtile_0__pin_dest_in_10_, right_width_0_height_3_subtile_0__pin_dest_in_11_, bottom_width_0_height_0_subtile_0__pin_dest_in_12_, bottom_width_0_height_0_subtile_0__pin_dest_in_13_, bottom_width_0_height_0_subtile_0__pin_dest_in_14_, bottom_width_0_height_0_subtile_0__pin_dest_in_15_, bottom_width_0_height_0_subtile_0__pin_dest_in_16_, bottom_width_0_height_0_subtile_0__pin_dest_in_17_, left_width_0_height_3_subtile_0__pin_dest_in_18_, left_width_0_height_3_subtile_0__pin_dest_in_19_, left_width_0_height_3_subtile_0__pin_dest_in_20_, left_width_0_height_3_subtile_0__pin_dest_in_21_, left_width_0_height_3_subtile_0__pin_dest_in_22_, left_width_0_height_3_subtile_0__pin_dest_in_23_}),
		.router_wrap_tile_is_tail_in({top_width_0_height_0_subtile_0__pin_is_tail_in_0_, bottom_width_0_height_0_subtile_0__pin_is_tail_in_1_, right_width_0_height_3_subtile_0__pin_is_tail_in_2_, left_width_0_height_3_subtile_0__pin_is_tail_in_3_}),
		.router_wrap_tile_send_in({top_width_0_height_0_subtile_0__pin_send_in_0_, bottom_width_0_height_0_subtile_0__pin_send_in_1_, right_width_0_height_3_subtile_0__pin_send_in_2_, left_width_0_height_3_subtile_0__pin_send_in_3_}),
		.router_wrap_tile_credit_in({top_width_0_height_0_subtile_0__pin_credit_in_0_, bottom_width_0_height_0_subtile_0__pin_credit_in_1_, right_width_0_height_3_subtile_0__pin_credit_in_2_, left_width_0_height_3_subtile_0__pin_credit_in_3_}),
		.router_wrap_tile_router_address({left_width_0_height_0_subtile_0__pin_router_address_0_, left_width_0_height_0_subtile_0__pin_router_address_1_, left_width_0_height_0_subtile_0__pin_router_address_2_, left_width_0_height_0_subtile_0__pin_router_address_3_}),
		.router_wrap_tile_axis_in_tvalid(left_width_0_height_1_subtile_0__pin_axis_in_tvalid_0_),
		.router_wrap_tile_axis_in_tdata({left_width_0_height_1_subtile_0__pin_axis_in_tdata_0_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_1_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_2_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_3_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_4_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_5_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_6_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_7_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_8_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_9_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_10_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_11_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_12_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_13_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_14_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_15_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_16_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_17_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_18_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_19_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_20_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_21_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_22_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_23_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_24_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_25_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_26_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_27_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_28_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_29_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_30_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_31_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_32_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_33_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_34_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_35_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_36_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_37_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_38_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_39_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_40_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_41_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_42_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_43_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_44_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_45_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_46_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_47_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_48_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_49_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_50_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_51_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_52_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_53_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_54_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_55_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_56_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_57_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_58_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_59_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_60_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_61_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_62_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_63_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_64_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_65_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_66_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_67_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_68_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_69_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_70_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_71_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_72_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_73_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_74_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_75_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_76_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_77_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_78_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_79_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_80_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_81_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_82_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_83_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_84_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_85_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_86_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_87_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_88_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_89_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_90_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_91_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_92_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_93_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_94_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_95_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_96_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_97_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_98_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_99_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_100_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_101_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_102_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_103_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_104_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_105_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_106_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_107_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_108_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_109_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_110_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_111_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_112_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_113_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_114_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_115_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_116_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_117_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_118_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_119_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_120_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_121_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_122_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_123_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_124_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_125_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_126_, left_width_0_height_1_subtile_0__pin_axis_in_tdata_127_}),
		.router_wrap_tile_axis_in_tlast(left_width_0_height_1_subtile_0__pin_axis_in_tlast_0_),
		.router_wrap_tile_axis_in_tid({left_width_0_height_1_subtile_0__pin_axis_in_tid_0_, left_width_0_height_1_subtile_0__pin_axis_in_tid_1_}),
		.router_wrap_tile_axis_in_tdest({right_width_0_height_1_subtile_0__pin_axis_in_tdest_0_, right_width_0_height_1_subtile_0__pin_axis_in_tdest_1_, right_width_0_height_1_subtile_0__pin_axis_in_tdest_2_, right_width_0_height_1_subtile_0__pin_axis_in_tdest_3_}),
		.router_wrap_tile_axis_out_tready(right_width_0_height_1_subtile_0__pin_axis_out_tready_0_),
		.router_wrap_tile_clk_usr(left_width_0_height_0_subtile_0__pin_clk_usr_0_),
		.ccff_head(ccff_head),
		.router_wrap_tile_credit_out({top_width_0_height_0_subtile_0__pin_credit_out_0_, bottom_width_0_height_0_subtile_0__pin_credit_out_1_, right_width_0_height_3_subtile_0__pin_credit_out_2_, left_width_0_height_3_subtile_0__pin_credit_out_3_}),
		.router_wrap_tile_data_out({top_width_0_height_0_subtile_0__pin_data_out_0_, top_width_0_height_0_subtile_0__pin_data_out_1_, top_width_0_height_0_subtile_0__pin_data_out_2_, top_width_0_height_0_subtile_0__pin_data_out_3_, top_width_0_height_0_subtile_0__pin_data_out_4_, top_width_0_height_0_subtile_0__pin_data_out_5_, top_width_0_height_0_subtile_0__pin_data_out_6_, top_width_0_height_0_subtile_0__pin_data_out_7_, top_width_0_height_0_subtile_0__pin_data_out_8_, top_width_0_height_0_subtile_0__pin_data_out_9_, top_width_0_height_0_subtile_0__pin_data_out_10_, top_width_0_height_0_subtile_0__pin_data_out_11_, top_width_0_height_0_subtile_0__pin_data_out_12_, top_width_0_height_0_subtile_0__pin_data_out_13_, top_width_0_height_0_subtile_0__pin_data_out_14_, top_width_0_height_0_subtile_0__pin_data_out_15_, top_width_0_height_0_subtile_0__pin_data_out_16_, top_width_0_height_0_subtile_0__pin_data_out_17_, top_width_0_height_0_subtile_0__pin_data_out_18_, top_width_0_height_0_subtile_0__pin_data_out_19_, top_width_0_height_0_subtile_0__pin_data_out_20_, top_width_0_height_0_subtile_0__pin_data_out_21_, top_width_0_height_0_subtile_0__pin_data_out_22_, top_width_0_height_0_subtile_0__pin_data_out_23_, top_width_0_height_0_subtile_0__pin_data_out_24_, top_width_0_height_0_subtile_0__pin_data_out_25_, top_width_0_height_0_subtile_0__pin_data_out_26_, top_width_0_height_0_subtile_0__pin_data_out_27_, top_width_0_height_0_subtile_0__pin_data_out_28_, top_width_0_height_0_subtile_0__pin_data_out_29_, top_width_0_height_0_subtile_0__pin_data_out_30_, top_width_0_height_0_subtile_0__pin_data_out_31_, bottom_width_0_height_0_subtile_0__pin_data_out_32_, bottom_width_0_height_0_subtile_0__pin_data_out_33_, bottom_width_0_height_0_subtile_0__pin_data_out_34_, bottom_width_0_height_0_subtile_0__pin_data_out_35_, bottom_width_0_height_0_subtile_0__pin_data_out_36_, bottom_width_0_height_0_subtile_0__pin_data_out_37_, bottom_width_0_height_0_subtile_0__pin_data_out_38_, bottom_width_0_height_0_subtile_0__pin_data_out_39_, bottom_width_0_height_0_subtile_0__pin_data_out_40_, bottom_width_0_height_0_subtile_0__pin_data_out_41_, bottom_width_0_height_0_subtile_0__pin_data_out_42_, bottom_width_0_height_0_subtile_0__pin_data_out_43_, bottom_width_0_height_0_subtile_0__pin_data_out_44_, bottom_width_0_height_0_subtile_0__pin_data_out_45_, bottom_width_0_height_0_subtile_0__pin_data_out_46_, bottom_width_0_height_0_subtile_0__pin_data_out_47_, bottom_width_0_height_0_subtile_0__pin_data_out_48_, bottom_width_0_height_0_subtile_0__pin_data_out_49_, bottom_width_0_height_0_subtile_0__pin_data_out_50_, bottom_width_0_height_0_subtile_0__pin_data_out_51_, bottom_width_0_height_0_subtile_0__pin_data_out_52_, bottom_width_0_height_0_subtile_0__pin_data_out_53_, bottom_width_0_height_0_subtile_0__pin_data_out_54_, bottom_width_0_height_0_subtile_0__pin_data_out_55_, bottom_width_0_height_0_subtile_0__pin_data_out_56_, bottom_width_0_height_0_subtile_0__pin_data_out_57_, bottom_width_0_height_0_subtile_0__pin_data_out_58_, bottom_width_0_height_0_subtile_0__pin_data_out_59_, bottom_width_0_height_0_subtile_0__pin_data_out_60_, bottom_width_0_height_0_subtile_0__pin_data_out_61_, bottom_width_0_height_0_subtile_0__pin_data_out_62_, bottom_width_0_height_0_subtile_0__pin_data_out_63_, right_width_0_height_3_subtile_0__pin_data_out_64_, right_width_0_height_3_subtile_0__pin_data_out_65_, right_width_0_height_3_subtile_0__pin_data_out_66_, right_width_0_height_3_subtile_0__pin_data_out_67_, right_width_0_height_3_subtile_0__pin_data_out_68_, right_width_0_height_3_subtile_0__pin_data_out_69_, right_width_0_height_3_subtile_0__pin_data_out_70_, right_width_0_height_3_subtile_0__pin_data_out_71_, right_width_0_height_3_subtile_0__pin_data_out_72_, right_width_0_height_3_subtile_0__pin_data_out_73_, right_width_0_height_3_subtile_0__pin_data_out_74_, right_width_0_height_3_subtile_0__pin_data_out_75_, right_width_0_height_3_subtile_0__pin_data_out_76_, right_width_0_height_3_subtile_0__pin_data_out_77_, right_width_0_height_3_subtile_0__pin_data_out_78_, right_width_0_height_3_subtile_0__pin_data_out_79_, right_width_0_height_3_subtile_0__pin_data_out_80_, right_width_0_height_3_subtile_0__pin_data_out_81_, right_width_0_height_3_subtile_0__pin_data_out_82_, right_width_0_height_3_subtile_0__pin_data_out_83_, right_width_0_height_3_subtile_0__pin_data_out_84_, right_width_0_height_3_subtile_0__pin_data_out_85_, right_width_0_height_3_subtile_0__pin_data_out_86_, right_width_0_height_3_subtile_0__pin_data_out_87_, right_width_0_height_3_subtile_0__pin_data_out_88_, right_width_0_height_3_subtile_0__pin_data_out_89_, right_width_0_height_3_subtile_0__pin_data_out_90_, right_width_0_height_3_subtile_0__pin_data_out_91_, right_width_0_height_3_subtile_0__pin_data_out_92_, right_width_0_height_3_subtile_0__pin_data_out_93_, right_width_0_height_3_subtile_0__pin_data_out_94_, right_width_0_height_3_subtile_0__pin_data_out_95_, left_width_0_height_3_subtile_0__pin_data_out_96_, left_width_0_height_3_subtile_0__pin_data_out_97_, left_width_0_height_3_subtile_0__pin_data_out_98_, left_width_0_height_3_subtile_0__pin_data_out_99_, left_width_0_height_3_subtile_0__pin_data_out_100_, left_width_0_height_3_subtile_0__pin_data_out_101_, left_width_0_height_3_subtile_0__pin_data_out_102_, left_width_0_height_3_subtile_0__pin_data_out_103_, left_width_0_height_3_subtile_0__pin_data_out_104_, left_width_0_height_3_subtile_0__pin_data_out_105_, left_width_0_height_3_subtile_0__pin_data_out_106_, left_width_0_height_3_subtile_0__pin_data_out_107_, left_width_0_height_3_subtile_0__pin_data_out_108_, left_width_0_height_3_subtile_0__pin_data_out_109_, left_width_0_height_3_subtile_0__pin_data_out_110_, left_width_0_height_3_subtile_0__pin_data_out_111_, left_width_0_height_3_subtile_0__pin_data_out_112_, left_width_0_height_3_subtile_0__pin_data_out_113_, left_width_0_height_3_subtile_0__pin_data_out_114_, left_width_0_height_3_subtile_0__pin_data_out_115_, left_width_0_height_3_subtile_0__pin_data_out_116_, left_width_0_height_3_subtile_0__pin_data_out_117_, left_width_0_height_3_subtile_0__pin_data_out_118_, left_width_0_height_3_subtile_0__pin_data_out_119_, left_width_0_height_3_subtile_0__pin_data_out_120_, left_width_0_height_3_subtile_0__pin_data_out_121_, left_width_0_height_3_subtile_0__pin_data_out_122_, left_width_0_height_3_subtile_0__pin_data_out_123_, left_width_0_height_3_subtile_0__pin_data_out_124_, left_width_0_height_3_subtile_0__pin_data_out_125_, left_width_0_height_3_subtile_0__pin_data_out_126_, left_width_0_height_3_subtile_0__pin_data_out_127_}),
		.router_wrap_tile_dest_out({top_width_0_height_0_subtile_0__pin_dest_out_0_, top_width_0_height_0_subtile_0__pin_dest_out_1_, top_width_0_height_0_subtile_0__pin_dest_out_2_, top_width_0_height_0_subtile_0__pin_dest_out_3_, top_width_0_height_0_subtile_0__pin_dest_out_4_, top_width_0_height_0_subtile_0__pin_dest_out_5_, right_width_0_height_3_subtile_0__pin_dest_out_6_, right_width_0_height_3_subtile_0__pin_dest_out_7_, right_width_0_height_3_subtile_0__pin_dest_out_8_, right_width_0_height_3_subtile_0__pin_dest_out_9_, right_width_0_height_3_subtile_0__pin_dest_out_10_, right_width_0_height_3_subtile_0__pin_dest_out_11_, bottom_width_0_height_0_subtile_0__pin_dest_out_12_, logical_tile_router_wrap_tile_mode_router_wrap_tile__0_undriven_router_wrap_tile_dest_out[13:17], left_width_0_height_3_subtile_0__pin_dest_out_18_, left_width_0_height_3_subtile_0__pin_dest_out_19_, left_width_0_height_3_subtile_0__pin_dest_out_20_, left_width_0_height_3_subtile_0__pin_dest_out_21_, left_width_0_height_3_subtile_0__pin_dest_out_22_, left_width_0_height_3_subtile_0__pin_dest_out_23_}),
		.router_wrap_tile_is_tail_out({top_width_0_height_0_subtile_0__pin_is_tail_out_0_, bottom_width_0_height_0_subtile_0__pin_is_tail_out_1_, right_width_0_height_3_subtile_0__pin_is_tail_out_2_, left_width_0_height_3_subtile_0__pin_is_tail_out_3_}),
		.router_wrap_tile_send_out({top_width_0_height_0_subtile_0__pin_send_out_0_, bottom_width_0_height_0_subtile_0__pin_send_out_1_, right_width_0_height_3_subtile_0__pin_send_out_2_, left_width_0_height_3_subtile_0__pin_send_out_3_}),
		.router_wrap_tile_axis_in_tready(right_width_0_height_0_subtile_0__pin_axis_in_tready_0_),
		.router_wrap_tile_axis_out_tvalid(right_width_0_height_1_subtile_0__pin_axis_out_tvalid_0_),
		.router_wrap_tile_axis_out_tdata({right_width_0_height_1_subtile_0__pin_axis_out_tdata_0_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_1_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_2_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_3_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_4_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_5_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_6_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_7_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_8_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_9_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_10_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_11_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_12_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_13_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_14_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_15_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_16_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_17_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_18_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_19_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_20_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_21_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_22_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_23_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_24_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_25_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_26_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_27_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_28_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_29_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_30_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_31_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_32_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_33_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_34_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_35_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_36_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_37_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_38_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_39_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_40_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_41_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_42_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_43_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_44_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_45_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_46_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_47_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_48_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_49_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_50_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_51_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_52_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_53_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_54_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_55_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_56_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_57_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_58_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_59_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_60_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_61_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_62_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_63_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_64_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_65_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_66_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_67_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_68_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_69_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_70_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_71_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_72_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_73_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_74_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_75_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_76_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_77_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_78_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_79_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_80_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_81_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_82_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_83_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_84_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_85_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_86_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_87_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_88_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_89_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_90_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_91_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_92_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_93_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_94_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_95_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_96_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_97_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_98_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_99_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_100_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_101_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_102_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_103_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_104_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_105_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_106_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_107_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_108_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_109_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_110_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_111_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_112_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_113_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_114_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_115_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_116_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_117_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_118_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_119_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_120_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_121_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_122_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_123_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_124_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_125_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_126_, right_width_0_height_1_subtile_0__pin_axis_out_tdata_127_}),
		.router_wrap_tile_axis_out_tlast(right_width_0_height_0_subtile_0__pin_axis_out_tlast_0_),
		.router_wrap_tile_axis_out_tid({right_width_0_height_0_subtile_0__pin_axis_out_tid_0_, right_width_0_height_0_subtile_0__pin_axis_out_tid_1_}),
		.router_wrap_tile_axis_out_tdest({right_width_0_height_0_subtile_0__pin_axis_out_tdest_0_, right_width_0_height_0_subtile_0__pin_axis_out_tdest_1_, right_width_0_height_0_subtile_0__pin_axis_out_tdest_2_, right_width_0_height_0_subtile_0__pin_axis_out_tdest_3_}),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_router_wrap_tile -----

//----- Default net type -----
`default_nettype wire



// ----- END Grid Verilog module: grid_router_wrap_tile -----

